`timescale 1ns/100ps

module adder(
);
	
endmodule
