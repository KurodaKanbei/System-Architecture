`timescale 100ns / 10ps

module loadRS (
	
);

endmodule
